module tb_quantizer();


   quantizer DUT(.*);
   
   initial begin
      
   end
endmodule // tb_quantizer
